
module test;







/*
    reg [3:0] mem [7:0]; // 8 x 4-bit vectors
    // reg [WIDTH-1:0] mem [DEPTH-1:0];


    initial begin
        for (int i=0; i<8; i++) begin
            mem[i] <= 0;
        end
    end

    always@(posedge clk or negedge res_n) begin
        if (~res_n) begin
            mem[i] <= 0;
        end else begin

        end
    end
*/
endmodule
